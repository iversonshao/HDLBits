module top_module( 
    input in, 
    output out 
);
//wire green;
//assign green = in;
assign out = in;

endmodule